magic
tech sky130A
timestamp 1720240049
<< nwell >>
rect -120 -120 120 225
<< nmos >>
rect -10 -300 5 -200
<< pmos >>
rect -10 -100 5 100
<< ndiff >>
rect -55 -210 -10 -200
rect -55 -290 -45 -210
rect -25 -290 -10 -210
rect -55 -300 -10 -290
rect 5 -210 50 -200
rect 5 -290 20 -210
rect 40 -290 50 -210
rect 5 -300 50 -290
<< pdiff >>
rect -45 90 -10 100
rect -45 -90 -40 90
rect -20 -90 -10 90
rect -45 -100 -10 -90
rect 5 90 40 100
rect 5 -90 15 90
rect 35 -90 40 90
rect 5 -100 40 -90
<< ndiffc >>
rect -45 -290 -25 -210
rect 20 -290 40 -210
<< pdiffc >>
rect -40 -90 -20 90
rect 15 -90 35 90
<< psubdiff >>
rect -60 -355 55 -340
rect -60 -390 -45 -355
rect 40 -390 55 -355
rect -60 -405 55 -390
<< nsubdiff >>
rect -55 190 50 200
rect -55 170 -40 190
rect 35 170 50 190
rect -55 160 50 170
<< psubdiffcont >>
rect -45 -390 40 -355
<< nsubdiffcont >>
rect -40 170 35 190
<< poly >>
rect -10 100 5 145
rect -10 -135 5 -100
rect -50 -145 5 -135
rect -50 -170 -40 -145
rect -15 -170 5 -145
rect -50 -180 5 -170
rect 60 -145 100 -135
rect 60 -170 70 -145
rect 95 -170 100 -145
rect 60 -180 100 -170
rect -10 -200 5 -180
rect -10 -325 5 -300
<< polycont >>
rect -40 -170 -15 -145
rect 70 -170 95 -145
<< locali >>
rect -55 195 50 200
rect -55 190 -25 195
rect 20 190 50 195
rect -55 170 -40 190
rect 35 170 50 190
rect -55 165 -25 170
rect 20 165 50 170
rect -55 160 50 165
rect -45 100 -20 160
rect -45 90 -15 100
rect -45 -90 -40 90
rect -20 -90 -15 90
rect -45 -100 -15 -90
rect 10 90 40 100
rect 10 -90 15 90
rect 35 -90 40 90
rect 10 -135 40 -90
rect -50 -145 -10 -135
rect -50 -170 -40 -145
rect -15 -170 -10 -145
rect -50 -180 -10 -170
rect 10 -145 100 -135
rect 10 -170 70 -145
rect 95 -170 100 -145
rect 10 -180 100 -170
rect 10 -200 40 -180
rect -55 -210 -15 -200
rect -55 -290 -45 -210
rect -25 -290 -15 -210
rect -55 -300 -15 -290
rect 10 -210 50 -200
rect 10 -290 20 -210
rect 40 -290 50 -210
rect 10 -300 50 -290
rect -55 -345 -25 -300
rect -55 -350 50 -345
rect -55 -355 -20 -350
rect 15 -355 50 -350
rect -55 -390 -45 -355
rect 40 -390 50 -355
rect -55 -395 -20 -390
rect 15 -395 50 -390
rect -55 -400 50 -395
rect -55 -405 -25 -400
<< viali >>
rect -25 190 20 195
rect -25 170 20 190
rect -25 165 20 170
rect -40 -170 -15 -145
rect 70 -170 95 -145
rect -20 -355 15 -350
rect -20 -390 15 -355
rect -20 -395 15 -390
<< metal1 >>
rect -320 195 310 200
rect -320 165 -25 195
rect 20 165 310 195
rect -320 160 310 165
rect -170 -145 0 -135
rect -170 -170 -40 -145
rect -15 -170 0 -145
rect -170 -180 0 -170
rect 15 -145 240 -135
rect 15 -170 70 -145
rect 95 -170 240 -145
rect 15 -180 240 -170
rect -305 -350 305 -340
rect -305 -395 -20 -350
rect 15 -395 305 -350
rect -305 -405 305 -395
<< labels >>
rlabel metal1 220 180 220 180 1 vdd
rlabel metal1 215 -160 220 -160 1 out
rlabel metal1 -145 -160 -140 -160 1 in
rlabel metal1 200 -375 205 -375 1 vss
<< end >>
